--RV32I_single Controls
--This is the controls for the RV32I_single design of the processor.
library IEEE;
 use IEEE.STD_LOGIC_1164.ALL;
 use IEEE.NUMERIC_STD.ALL;
entity RV32I_single is
Port(
	--Error Signal
		error: out std_logic;	--Instruction
		instr: in std_logic_vector(31 downto 0);

	--Control Signals
		mux_reg_write : out std_logic_vector(1 downto 0);
		mux_output : out std_logic;
		mux_reg_descr_alu : out std_logic;
		mux_reg_pc_alu : out std_logic;
		control_mem_writeenable : out std_logic;
		control_alu : out std_logic_vector(3 downto 0);
		control_reg_writeenable : out std_logic;
		control_branch : out std_logic_vector(3 downto 0);
		control_mem_logic : out std_logic_vector(3 downto 0));
end RV32I_single;
architecture Controls_Behavior of RV32I_single is


begin
	RV32I_single_process : process(instr)
		begin
				case instr(6 downto 0)&instr(14 downto 12)&instr(30) is
					when "00000110000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0000";
						error <= '0';
					when "00000110001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0000";
						error <= '0';
					when "00000110010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0001";
						error <= '0';
					when "00000110011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0001";
						error <= '0';
					when "00000110100" =>
						mux_reg_write <= "00";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0010";
						error <= '0';
					when "00000110101" =>
						mux_reg_write <= "00";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0010";
						error <= '0';
					when "00000111000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0100";
						error <= '0';
					when "00000111001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0100";
						error <= '0';
					when "00000111010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0101";
						error <= '0';
					when "00000111011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "0101";
						error <= '0';
					when "00011110000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00011110001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00011110010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00011110011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110001" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0001";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0010";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110101" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0010";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0011";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100110111" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0011";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0100";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111001" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0100";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0101";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111011" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1101";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0110";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111101" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0110";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0111";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00100111111" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0111";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110001" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110011" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110101" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101110111" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111001" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111011" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111101" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "00101111111" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01000110000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1000";
						error <= '0';
					when "01000110001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1000";
						error <= '0';
					when "01000110010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1001";
						error <= '0';
					when "01000110011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1001";
						error <= '0';
					when "01000110100" =>
						mux_reg_write <= "00";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1010";
						error <= '0';
					when "01000110101" =>
						mux_reg_write <= "00";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '1';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1010";
						error <= '0';
					when "01100110000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100110001" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100110010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0001";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100110100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0010";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100110110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0011";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100111000" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0100";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100111010" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0101";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100111011" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "1101";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100111100" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0110";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01100111110" =>
						mux_reg_write <= "11";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0111";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110000" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110001" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110010" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110011" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110100" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110101" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110110" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101110111" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111000" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111001" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111010" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111011" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111100" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111101" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111110" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "01101111111" =>
						mux_reg_write <= "11";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000110000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1000";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000110001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1000";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000110010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1001";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000110011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1001";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1100";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1100";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1101";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1101";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111100" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1110";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111101" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1110";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111110" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1111";
						control_mem_logic <= "1111";
						error <= '0';
					when "11000111111" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "1000";
						control_reg_writeenable <= '0';
						control_branch <= "1111";
						control_mem_logic <= "1111";
						error <= '0';
					when "11001110000" =>
						mux_reg_write <= "01";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0001";
						control_mem_logic <= "1111";
						error <= '0';
					when "11001110001" =>
						mux_reg_write <= "01";
						mux_output <= '0';
						mux_reg_descr_alu <= '1';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0001";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110000" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110001" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110010" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110011" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110100" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110101" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110110" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011110111" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111000" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111001" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111010" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111011" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111100" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111101" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111110" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11011111111" =>
						mux_reg_write <= "01";
						mux_output <= '1';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '1';
						control_branch <= "0011";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110000" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110001" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110100" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110101" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110110" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100110111" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111010" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111011" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111100" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111101" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111110" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when "11100111111" =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '0';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '0';
					when others =>
						mux_reg_write <= "10";
						mux_output <= '0';
						mux_reg_descr_alu <= '0';
						mux_reg_pc_alu <= '1';
						control_mem_writeenable <= '0';
						control_alu <= "0000";
						control_reg_writeenable <= '0';
						control_branch <= "0010";
						control_mem_logic <= "1111";
						error <= '1';
				end case;
	end process RV32I_single_process;
end Controls_Behavior;
